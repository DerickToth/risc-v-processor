module risc_processor(clk);
endmodule