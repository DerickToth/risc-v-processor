module risc_processor(clk50);
	
	wire clk80
	
	
	always @(*): begin
		//combinational logic blocks
	end
	
	always@(posedge clk80): begin
		//x = next_x
	end
	
	always@(negedge clk80): begin
		//x = next_x
	end
endmodule