module immediateGenerator();
endmodule