module registerFile();
endmodule